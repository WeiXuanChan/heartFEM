*version 4.0.0
*units in Pressure:mmHg, Volume:mL, time:ms
*chamber source mode: 0=pressure pulse with capacitor, 1=fourier current, 2=timebased, 3=2d table,4=2dtable with trackphase, 5=3d table ,6=3dtable with trackphase
.title LV full circuit

.PARAM PI = 3.14159265359
.PARAM lasourcemode = <<lasourcemode>>
.PARAM rasourcemode = <<rasourcemode>>
.PARAM lvsourcemode = <<lvsourcemode>>
.PARAM rvsourcemode = <<rvsourcemode>>

.func manmod(shorttime,period) {shorttime - floor(shorttime / period) * period}
.func disfrompeak(xtime,peaktime,width,period) {min( abs( xtime - peaktime) , period - abs( xtime - peaktime))}
.func cossq(xtime,amp,peaktime,width,period) {amp * cos( PI * disfrompeak( xtime , peaktime , width,period ) / width)^2}

.model valve sidiode(Roff=10meg Ron=1 Rrev=10k Vfwd=0.1 Vrev=1k Revepsilon=0.2 Epsilon=0.2)

.subckt vein in out rval=100meg lval=1m
R1 1  out    r = rval
L1 in 1    l = lval
.ends vein

Eheartperiod heartperiod gnd vol = ' <<cycle>> '
Bcumulativeheartphase  cumulativeheartphase gnd I = -2*PI/v(heartperiod) 
acumulativeheartphase  cumulativeheartphase gnd heartphaseconvertcap
.model heartphaseconvertcap capacitor (c=1 ic=0)
Eheartphase heartphase gnd vol = ' manmod(v(cumulativeheartphase),2*PI) '
Elaactivepeaktime laactivepeaktime gnd vol = ' <<latimetopeaktension>> '
Eraactivepeaktime raactivepeaktime gnd vol = ' <<ratimetopeaktension>> '
Elvactivepeaktime lvactivepeaktime gnd vol = ' <<lvtimetopeaktension>> '
Ervactivepeaktime rvactivepeaktime gnd vol = ' <<rvtimetopeaktension>> '
Elvregurgitationvalveratio lvregurgitationvalveratio gnd vol = ' <<lvregurgevalveratio>> '
Eaaregurgitationvalveratio aaregurgitationvalveratio gnd vol = ' <<aaregurgevalveratio>> '
Ervregurgitationvalveratio rvregurgitationvalveratio gnd vol = ' <<rvregurgevalveratio>> '
Epa1regurgitationvalveratio pa1regurgitationvalveratio gnd vol = ' <<pa1regurgevalveratio>> '
Etime timecyclic gnd vol = 'v(heartperiod) *v(heartphase)/2/PI'

Vlaprobe la    lagnd  dc 0
Vraprobe ra    ragnd dc 0
Vlvprobe lv    lvgnd  dc 0
Vrvprobe rv    rvgnd dc 0

.if (lasourcemode == 0)
Cla    lagnd   lagnd2   <<lac>> 
Elau   lagnd2  gnd      vol = 'cossq( v(timecyclic) ,<<laamp>>,<<lapeaktime>>,<<lawidth>>,v(heartperiod))'
Vpasslaphasetime laphasetime timecyclic dc 0
.elseif (lasourcemode == 1)
Glau1   lagnd       gnd   cur = '<<lauamp1>> * sin(manmod(v(cumulativeheartphase),2*PI) +       <<lauphase1>>/180*PI)'
Glau2   lagnd       gnd   cur = '<<lauamp2>> * sin(manmod(v(cumulativeheartphase),PI) * 2 +     <<lauphase2>>/180*PI)'
Glau3   lagnd       gnd   cur = '<<lauamp3>> * sin(manmod(v(cumulativeheartphase),PI*2/3) * 3 + <<lauphase3>>/180*PI)'
Glau4   lagnd       gnd   cur = '<<lauamp4>> * sin(manmod(v(cumulativeheartphase),PI/2) * 4 +   <<lauphase4>>/180*PI)'
Vpasslaphasetime laphasetime timecyclic dc 0
.else
Blau   lagnd   gnd  <<lainputvar>> = v(lagenerator0) + v(lagenerator1)
.if (lasourcemode == 2)
alau0 %v[lagenerator0] la_pwl_input
.model la_pwl_input filesource (file="<<laufile>>" amploffset=[0] amplscale=[1] timeoffset=0 timescale=1 timerelative=false amplstep=false)
Vlau1 lagenerator1   gnd  dc 0
Vpasslaphasetime laphasetime timecyclic dc 0
.else
.if (lasourcemode < 5)
alau0 gnd lavol %v(lagenerator0) lautabmod0
.model lautabmod0 table2d (offset=0.0 gain=1 order=3 file="<<lautablebasefile>>")
alau1 lavol laphasetime %v(lagenerator1) lautabmod
.model lautabmod table2d (offset=0.0 gain=1 order=3 file="<<lautablefile>>")
.else
alau0 ravol lavol %v(lagenerator0) lautabmod0
.model lautabmod0 table2d (offset=0.0 gain=1 order=3 file="<<lautablebasefile>>")
alau1 lavol laphasetime ravol %v(lagenerator1) lautabmod
.model lautabmod table3d (offset=0.0 gain=1 order=3 file="<<lautablefile>>")
.endif
.if (lasourcemode == 3 || lasourcemode == 5)
Vpasslaphasetime laphasetime timecyclic dc 0
.else
Bestphase laestphase gnd V = v(timecyclic)/v(laactivepeaktime)
Blarisecurrent gnd lacurrentphase I =  ((v(timecyclic) <= v(laactivepeaktime)) ? (v(lacurrentphase) >= (1 - (3 * <<stepTime>> * v(larisetemp)))  ? (1-v(lacurrentphase))/(3 * <<stepTime>> * v(larisetemp))*v(larisetemp) : v(larisetemp) ) : 0)
Blarisetemp larisetemp gnd V = 1/v(laactivepeaktime)*10
Blafallcurrent lacurrentphase gnd I = (v(timecyclic) < v(laactivepeaktime)) ? 0 : v(lafalltemp)
Blafalltemp lafalltemp gnd V =  1/v(latr)
alapressgrad  lacurrentphase gnd latrcap
.model latrcap capacitor (c=1 ic=0)
.if (lasourcemode == 4)
alatr gnd lavol %v(latr) lautabtrmod
.model lautabtrmod table2d (offset=0.0 gain=1 order=3 file="<<latrtablefile>>")
.else
alatr ravol lavol %v(latr) lautabtrmod
.model lautabtrmod table2d (offset=0.0 gain=1 order=3 file="<<latrtablefile>>")
.endif
Blaphase laphase gnd V = max(0,min(1,v(lacurrentphase)))
Btime2 laphasetime gnd V =  (v(timecyclic) > v(laactivepeaktime)) ? (v(laactivepeaktime) + v(latr) * (1-v(lacurrentphase))) : v(timecyclic)
.endif
.endif
.endif


.if (rasourcemode == 0)
Cra    ragnd   ragnd2   <<rac>> 
Erau   ragnd2  gnd      vol = 'cossq( v(timecyclic) ,<<raamp>>,<<rapeaktime>>,<<rawidth>>,v(heartperiod))'
Vpassraphasetime raphasetime timecyclic dc 0
.elseif (rasourcemode == 1)
Grau1   ragnd       gnd   cur = '<<rauamp1>> * sin(manmod(v(cumulativeheartphase),2*PI) +       <<rauphase1>>/180*PI)'
Grau2   ragnd       gnd   cur = '<<rauamp2>> * sin(manmod(v(cumulativeheartphase),PI) * 2 +     <<rauphase2>>/180*PI)'
Grau3   ragnd       gnd   cur = '<<rauamp3>> * sin(manmod(v(cumulativeheartphase),PI*2/3) * 3 + <<rauphase3>>/180*PI)'
Grau4   ragnd       gnd   cur = '<<rauamp4>> * sin(manmod(v(cumulativeheartphase),PI/2) * 4 +   <<rauphase4>>/180*PI)'
Vpassraphasetime raphasetime timecyclic dc 0
.else
Brau   ragnd   gnd  <<rainputvar>> = v(ragenerator0) + v(ragenerator1)
.if (rasourcemode == 2)
arau0 %v[ragenerator0] ra_pwl_input
.model ra_pwl_input filesource (file="<<raufile>>" amploffset=[0] amplscale=[1] timeoffset=0 timescale=1 timerelative=false amplstep=false)
Vrau1 ragenerator1   gnd  dc 0
Vpassraphasetime raphasetime timecyclic dc 0
.else
.if (rasourcemode < 5)
arau0 gnd ravol %v(ragenerator0) rautabmod0
.model rautabmod0 table2d (offset=0.0 gain=1 order=3 file="<<rautablebasefile>>")
arau1 ravol raphasetime %v(ragenerator1) rautabmod
.model rautabmod table2d (offset=0.0 gain=1 order=3 file="<<rautablefile>>")
.else
arau0 ravol lavol %v(ragenerator0) rautabmod0
.model rautabmod0 table2d (offset=0.0 gain=1 order=3 file="<<rautablebasefile>>")
arau1 lavol raphasetime ravol %v(ragenerator1) rautabmod
.model rautabmod table3d (offset=0.0 gain=1 order=3 file="<<rautablefile>>")
.endif
.if (rasourcemode == 3 || rasourcemode == 5)
Vpassraphasetime raphasetime timecyclic dc 0
.else
Bestphase raestphase gnd V = v(timecyclic)/v(raactivepeaktime)
Brarisecurrent gnd racurrentphase I =  ((v(timecyclic) <= v(raactivepeaktime)) ? (v(racurrentphase) >= (1 - (3 * <<stepTime>> * v(rarisetemp)))  ? (1-v(racurrentphase))/(3 * <<stepTime>> * v(rarisetemp))*v(rarisetemp) : v(rarisetemp) ) : 0)
Brarisetemp rarisetemp gnd V = 1/v(raactivepeaktime)*10
Brafallcurrent racurrentphase gnd I = (v(timecyclic) < v(raactivepeaktime)) ? 0 : v(rafalltemp)
Brafalltemp rafalltemp gnd V =  1/v(ratr)
arapressgrad  racurrentphase gnd ratrcap
.model ratrcap capacitor (c=1 ic=0)
.if (rasourcemode == 4)
aratr gnd ravol %v(ratr) rautabtrmod
.model rautabtrmod table2d (offset=0.0 gain=1 order=3 file="<<ratrtablefile>>")
.else
aratr ravol lavol %v(ratr) rautabtrmod
.model rautabtrmod table2d (offset=0.0 gain=1 order=3 file="<<ratrtablefile>>")
.endif
Braphase raphase gnd V = max(0,min(1,v(racurrentphase)))
Btime2 raphasetime gnd V =  (v(timecyclic) > v(raactivepeaktime)) ? (v(raactivepeaktime) + v(ratr) * (1-v(racurrentphase))) : v(timecyclic)
.endif
.endif
.endif

.if (lvsourcemode == 0)
Clv    lvgnd   lvgnd2   <<lvc>> 
Elvu   lvgnd2  gnd      vol = 'cossq( v(timecyclic) ,<<lvamp>>,<<lvpeaktime>>,<<lvwidth>>,v(heartperiod))'
Vpasslvphasetime lvphasetime timecyclic dc 0
.elseif (lvsourcemode == 1)
Glvu1   lvgnd       gnd   cur = '<<lvuamp1>> * sin(manmod(v(cumulativeheartphase),2*PI) +       <<lvuphase1>>/180*PI)'
Glvu2   lvgnd       gnd   cur = '<<lvuamp2>> * sin(manmod(v(cumulativeheartphase),PI) * 2 +     <<lvuphase2>>/180*PI)'
Glvu3   lvgnd       gnd   cur = '<<lvuamp3>> * sin(manmod(v(cumulativeheartphase),PI*2/3) * 3 + <<lvuphase3>>/180*PI)'
Glvu4   lvgnd       gnd   cur = '<<lvuamp4>> * sin(manmod(v(cumulativeheartphase),PI/2) * 4 +   <<lvuphase4>>/180*PI)'
Vpasslvphasetime lvphasetime timecyclic dc 0
.else
Blvu   lvgnd   gnd  <<lvinputvar>> = v(lvgenerator0) + v(lvgenerator1)
.if (lvsourcemode == 2)
alvu0 %v[lvgenerator0] lv_pwl_input
.model lv_pwl_input filesource (file="<<lvufile>>" amploffset=[0] amplscale=[1] timeoffset=0 timescale=1 timerelative=false amplstep=false)
Vlvu1 lvgenerator1   gnd  dc 0
Vpasslvphasetime lvphasetime timecyclic dc 0
.else
.if (lvsourcemode < 5)
alvu0 gnd lvvol %v(lvgenerator0) lvutabmod0
.model lvutabmod0 table2d (offset=0.0 gain=1 order=3 file="<<lvutablebasefile>>")
alvu1 lvvol lvphasetime %v(lvgenerator1) lvutabmod
.model lvutabmod table2d (offset=0.0 gain=1 order=3 file="<<lvutablefile>>")
.else
alvu0 rvvol lvvol %v(lvgenerator0) lvutabmod0
.model lvutabmod0 table2d (offset=0.0 gain=1 order=3 file="<<lvutablebasefile>>")
alvu1 lvvol lvphasetime rvvol %v(lvgenerator1) lvutabmod
.model lvutabmod table3d (offset=0.0 gain=1 order=3 file="<<lvutablefile>>")
.endif
.if (lvsourcemode == 3 || lvsourcemode == 5)
Vpasslvphasetime lvphasetime timecyclic dc 0
.else
Bestphase lvestphase gnd V = v(timecyclic)/v(lvactivepeaktime)
Blvrisecurrent gnd lvcurrentphase I =  ((v(timecyclic) <= v(lvactivepeaktime)) ? (v(lvcurrentphase) >= (1 - (3 * <<stepTime>> * v(lvrisetemp)))  ? (1-v(lvcurrentphase))/(3 * <<stepTime>> * v(lvrisetemp))*v(lvrisetemp) : v(lvrisetemp) ) : 0)
Blvrisetemp lvrisetemp gnd V = 1/v(lvactivepeaktime)*10
Blvfallcurrent lvcurrentphase gnd I = (v(timecyclic) < v(lvactivepeaktime)) ? 0 : v(lvfalltemp)
Blvfalltemp lvfalltemp gnd V =  1/v(lvtr)
alvpressgrad  lvcurrentphase gnd lvtrcap
.model lvtrcap capacitor (c=1 ic=0)
.if (lvsourcemode == 4)
alvtr gnd lvvol %v(lvtr) lvutabtrmod
.model lvutabtrmod table2d (offset=0.0 gain=1 order=3 file="<<lvtrtablefile>>")
.else
alvtr rvvol lvvol %v(lvtr) lvutabtrmod
.model lvutabtrmod table2d (offset=0.0 gain=1 order=3 file="<<lvtrtablefile>>")
.endif
Blvphase lvphase gnd V = max(0,min(1,v(lvcurrentphase)))
Btime2 lvphasetime gnd V =  (v(timecyclic) > v(lvactivepeaktime)) ? (v(lvactivepeaktime) + v(lvtr) * (1-v(lvcurrentphase))) : v(timecyclic)
.endif
.endif
.endif

.if (rvsourcemode == 0)
Crv    rvgnd   rvgnd2   <<rvc>> 
Ervu   rvgnd2  gnd      vol = 'cossq( v(timecyclic) ,<<rvamp>>,<<rvpeaktime>>,<<rvwidth>>,v(heartperiod))'
Vpassrvphasetime rvphasetime timecyclic dc 0
.elseif (rvsourcemode == 1)
Grvu1   rvgnd       gnd   cur = '<<rvuamp1>> * sin(manmod(v(cumulativeheartphase),2*PI) +       <<rvuphase1>>/180*PI)'
Grvu2   rvgnd       gnd   cur = '<<rvuamp2>> * sin(manmod(v(cumulativeheartphase),PI) * 2 +     <<rvuphase2>>/180*PI)'
Grvu3   rvgnd       gnd   cur = '<<rvuamp3>> * sin(manmod(v(cumulativeheartphase),PI*2/3) * 3 + <<rvuphase3>>/180*PI)'
Grvu4   rvgnd       gnd   cur = '<<rvuamp4>> * sin(manmod(v(cumulativeheartphase),PI/2) * 4 +   <<rvuphase4>>/180*PI)'
Vpassrvphasetime rvphasetime timecyclic dc 0
.else
Brvu   rvgnd   gnd  <<rvinputvar>> = v(rvgenerator0) + v(rvgenerator1)
.if (rvsourcemode == 2)
arvu0 %v[rvgenerator0] rv_pwl_input
.model rv_pwl_input filesource (file="<<rvufile>>" amploffset=[0] amplscale=[1] timeoffset=0 timescale=1 timerelative=false amplstep=false)
Vrvu1 rvgenerator1   gnd  dc 0
Vpassrvphasetime rvphasetime timecyclic dc 0
.else
.if (rvsourcemode <5)
arvu0 gnd rvvol %v(rvgenerator0) rvutabmod0
.model rvutabmod0 table2d (offset=0.0 gain=1 order=3 file="<<rvutablebasefile>>")
arvu1 rvvol rvphasetime %v(rvgenerator1) rvutabmod
.model rvutabmod table2d (offset=0.0 gain=1 order=3 file="<<rvutablefile>>")
.else
arvu0 rvvol lvvol %v(rvgenerator0) rvutabmod0
.model rvutabmod0 table2d (offset=0.0 gain=1 order=3 file="<<rvutablebasefile>>")
arvu1 lvvol rvphasetime rvvol %v(rvgenerator1) rvutabmod
.model rvutabmod table3d (offset=0.0 gain=1 order=3 file="<<rvutablefile>>")
.endif
.if (rvsourcemode == 3 || rvsourcemode == 5)
Vpassrvphasetime rvphasetime timecyclic dc 0
.else
Bestphase rvestphase gnd V = v(timecyclic)/v(rvactivepeaktime)
Brvrisecurrent gnd rvcurrentphase I =  ((v(timecyclic) <= v(rvactivepeaktime)) ? (v(rvcurrentphase) >= (1 - (3 * <<stepTime>> * v(rvrisetemp)))  ? (1-v(rvcurrentphase))/(3 * <<stepTime>> * v(rvrisetemp))*v(rvrisetemp) : v(rvrisetemp) ) : 0)
Brvrisetemp rvrisetemp gnd V = 1/v(rvactivepeaktime)*10
Brvfallcurrent rvcurrentphase gnd I = (v(timecyclic) < v(rvactivepeaktime)) ? 0 : v(rvfalltemp)
Brvfalltemp rvfalltemp gnd V =  1/v(rvtr)
arvpressgrad  rvcurrentphase gnd rvtrcap
.model rvtrcap capacitor (c=1 ic=0)
.if (rvsourcemode == 4)
arvtr gnd rvvol %v(rvtr) rvutabtrmod
.model rvutabtrmod table2d (offset=0.0 gain=1 order=3 file="<<rvtrtablefile>>")
.else
arvtr rvvol lvvol %v(rvtr) rvutabtrmod
.model rvutabtrmod table2d (offset=0.0 gain=1 order=3 file="<<rvtrtablefile>>")
.endif
Brvphase rvphase gnd V = max(0,min(1,v(rvcurrentphase)))
Btime2 rvphasetime gnd V =  (v(timecyclic) > v(rvactivepeaktime)) ? (v(rvactivepeaktime) + v(rvtr) * (1-v(rvcurrentphase))) : v(timecyclic)
.endif
.endif
.endif


Blavol  lavol gnd I = -i(Vlaprobe) 
alavolconvert  lavol gnd lavolconvertcap
.model lavolconvertcap capacitor (c=1 ic=<<lainitvol>>)

Bravol  ravol gnd I = -i(Vraprobe) 
aravolconvert  ravol gnd ravolconvertcap
.model ravolconvertcap capacitor (c=1 ic=<<rainitvol>>)

Blvvol  lvvol gnd I = -i(Vlvprobe) 
alvvolconvert  lvvol gnd lvvolconvertcap
.model lvvolconvertcap capacitor (c=1 ic=<<lvinitvol>>)

Brvvol  rvvol gnd I = -i(Vrvprobe) 
arvvolconvert  rvvol gnd rvvolconvertcap
.model rvvolconvertcap capacitor (c=1 ic=<<rvinitvol>>)

Vlalavalv  lavalvp1 lavalvp2 dc 0
Vlvlvvalv  lv  lvvalvp1 dc 0
Vraravalv  ravalvp1 ravalvp2 dc 0
Vrvrvvalv  rv  rvvalvp1 dc 0
Vfo  fovalvp1 fovalvp2 dc 0
Vda  ao2p1 ao2p2 dc 0
Vdv  ivcp1 ivcp2 dc 0

Elalavalvk lalavalvk gnd vol = ' <<lalavalvk>> '
Blalavalv  lavalvp2 lavalv V=' v(lalavalvk) * ( i(Vlalavalv) ^2 )^( <<lalavalvb>> / 2) * sgn( i(Vlalavalv) ) '
Elvlvvalvk lvlvvalvk gnd vol = ' <<lvlvvalvk>> '
Blvlvvalv  lvvalvp1 lvvalvp2 V=' v(lvlvvalvk) * ( i(Vlvlvvalv) ^2 )^( <<lvlvvalvb>> / 2) * sgn( i(Vlvlvvalv) ) '
Eraravalvk raravalvk gnd vol = ' <<raravalvk>> '
Braravalv  ravalvp2 ravalv V=' v(raravalvk) * ( i(Vraravalv) ^2 )^( <<raravalvb>> / 2) * sgn( i(Vraravalv) ) '
Ervrvvalvk rvrvvalvk gnd vol = ' <<rvrvvalvk>> '
Brvrvvalv  rvvalvp1 rvvalvp2 V=' v(rvrvvalvk) * ( i(Vrvrvvalv) ^2 )^( <<rvrvvalvb>> / 2) * sgn( i(Vrvrvvalv) ) '
Efok fok gnd vol = ' <<fok>> '
Bfo  fovalvp2 fovalv V=' v(fok) * ( i(Vfo) ^2 )^( <<fob>> / 2) * sgn( i(Vfo) ) '
Edak dak gnd vol = ' <<dak>> '
Bda  ao2p2 ao2 V=' v(dak) * ( i(Vda) ^2 )^( <<dab>> / 2) * sgn( i(Vda) ) '
Edvk dvk gnd vol = ' <<dvk>> '
Bdv  ivcp2 ivc V=' v(dvk) * ( i(Vdv) ^2 )^( <<dvb>> / 2) * sgn( i(Vdv) ) '

ala   lavalv   lv      valve
alv   lvvalvp2 lvvalv  valve
ara   ravalv   rv    valve
arv   rvvalvp2 rvvalv    valve
afo   fovalv   la    valve


Vlvregurgitation  lv          lvregurp1   dc 0
Blvregurgitation  lvregurp1   lvregurp2   V=' v(lalavalvk) / max(v(lvregurgitationvalveratio),1n) * ( i(Vlvregurgitation) ^2 )^( <<lalavalvb>> / 2) * sgn( i(Vlvregurgitation) ) '
alvregurgitation  lvregurp2   lavalvp1    valve

Vaaregurgitation  lvvalv      aaregurp1   dc 0
Baaregurgitation  aaregurp1   aaregurp2   V=' v(lvlvvalvk) / max(v(aaregurgitationvalveratio),1n) * ( i(Vaaregurgitation) ^2 )^( <<lvlvvalvb>> / 2) * sgn( i(Vaaregurgitation) ) '
aaaregurgitation  aaregurp2   lv    valve

Vrvregurgitation  rv          rvregurp1   dc 0
Brvregurgitation  rvregurp1   rvregurp2   V=' v(raravalvk) / max(v(rvregurgitationvalveratio),1n) * ( i(Vrvregurgitation) ^2 )^( <<raravalvb>> / 2) * sgn( i(Vrvregurgitation) ) '
arvregurgitation  rvregurp2   ravalvp1    valve

Vpa1regurgitation  rvvalv       pa1regurp1   dc 0
Bpa1regurgitation  pa1regurp1   pa1regurp2   V=' v(rvrvvalvk) / max(v(pa1regurgitationvalveratio),1n) * ( i(Vpa1regurgitation) ^2 )^( <<rvrvvalvb>> / 2) * sgn( i(Vpa1regurgitation) ) '
apa1regurgitation  pa1regurp2   ravalvp1    valve


Caa   aa    gnd    <<aac>>    
Cao1  ao1   gnd    <<ao1c>>   
Cao2  ao2   gnd    <<ao2c>>   
Cao3  ao3   gnd    <<ao3c>>   
Cao4  ao4   gnd    <<ao4c>>   
Cbr   br    gnd    <<brc>>    
Cca   ca    gnd    <<cac>>    
Cub   ub    gnd    <<ubc>>    
Che   he    gnd    <<hec>>    
Cinte inte  gnd    <<intec>> 
Civc  ivc   gnd    <<ivcc>>   
Ckid  kid   gnd    <<kidc>>  
Cleg  leg   gnd    <<legc>>   
Clung lung  gnd    <<lungc>>  
Cpa1  pa1   gnd    <<pa1c>>   
Cpa2  pa2   gnd    <<pa2c>>   
Cplac plac  gnd    <<placc>>  
Csvc  svc   gnd    <<svcc>>  
Cuv   uv    gnd    <<uvc>>   

Xlalavalv  la  lavalvp1    vein  rval=<<lalavalvr>>    lval=<<lalavalvl>>
Xlvlvvalv  lvvalv   aa    vein  rval=<<lvlvvalvr>>    lval=<<lvlvvalvl>>
Xraravalv  ra  ravalvp1    vein  rval=<<raravalvr>>    lval=<<raravalvl>>
Xrvrvvalv  rvvalv   pa1   vein  rval=<<rvrvvalvr>>    lval=<<rvrvvalvl>>


Xcabr     ca    br     vein  rval=<<cabrr>>     lval=<<cabrl>>
Xbrsvc    br    svc    vein  rval=<<brsvcr>>    lval=<<brsvcl>>
Xubsvc    ub    svc    vein  rval=<<ubsvcr>>    lval=<<ubsvcl>>
Xao1ca    ao1   ca     vein  rval=<<ao1car>>    lval=<<ao1cal>>
Xao1ub    ao1   ub     vein  rval=<<ao1ubr>>    lval=<<ao1ubl>>
Xsvcra    svc   ra     vein  rval=<<svcrar>>    lval=<<svcral>>
Xpa1pa2   pa1   pa2    vein  rval=<<pa1pa2r>>   lval=<<pa1pa2l>>
Xpa2lung  pa2   lung   vein  rval=<<pa2lungr>>  lval=<<pa2lungl>>
Xlungla   lung  la     vein  rval=<<lunglar>>   lval=<<lunglal>>
Xaaao1    aa    ao1    vein  rval=<<aaao1r>>    lval=<<aaao1l>>
Xao1ao2   ao1   ao2    vein  rval=<<ao1ao2r>>   lval=<<ao1ao2l>>
Xao2ao3   ao2   ao3    vein  rval=<<ao2ao3r>>   lval=<<ao2ao3l>>
Xao3ao4   ao3   ao4    vein  rval=<<ao3ao4r>>   lval=<<ao3ao4l>>
Xao3kid   ao3   kid    vein  rval=<<ao3kidr>>   lval=<<ao3kidl>>
Xao3he    ao3   he     vein  rval=<<ao3her>>    lval=<<ao3hel>>
Xao3inte  ao3   inte   vein  rval=<<ao3inter>>  lval=<<ao3intel>>
Xao4leg   ao4   leg    vein  rval=<<ao4legr>>   lval=<<ao4legl>>
Xao4plac  ao4   plac   vein  rval=<<ao4placr>>  lval=<<ao4placl>>
Xkidivc   kid   ivc    vein  rval=<<kidivcr>>   lval=<<kidivcl>>
Xintehe   inte  he     vein  rval=<<inteher>>   lval=<<intehel>>
Xlegivc   leg   ivc    vein  rval=<<legivcr>>   lval=<<legivcl>>
Xplacuv   plac  uv     vein  rval=<<placuvr>>   lval=<<placuvl>>
Xuvhe     uv    he     vein  rval=<<uvher>>     lval=<<uvhel>>
Xheivc    he    ivc    vein  rval=<<heivcr>>    lval=<<heivcl>>
Xivcra    ivc   ra     vein  rval=<<ivcrar>>    lval=<<ivcral>>

Xda       pa2   ao2p1    vein  rval=<<dar>>    lval=<<dal>>
Xdv       uv    ivcp1    vein  rval=<<dvr>>    lval=<<dvl>>
Xfo       ivc   fovalvp1 vein  rval=<<for>>    lval=<<fol>>


.options savecurrents

.ic v(la)= <<vla0>> v(ra)= <<vra0>>
.tran <<stepTime>> <<stopTime>>
*.print tran v(lv) i(Vlvprobe)


.control
set controlswait
set filetype=ascii
set wr_vecnames
run
wrdata <<outfile>> v(lv) v(lvvol) v(la) v(rv) v(ra) v(pa1) v(aa) v(lavalvp1) v(lvvalv) i(Vlvprobe) v(lvphasetime) v(rvvol) i(Vlalavalv) i(Vlvlvvalv) i(Vlvregurgitation) v(lvregurp2) v(lvvalvp2) i(Vrvprobe)
.endc 
.end
