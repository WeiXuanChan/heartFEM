*version 3.1.2

.title LV full circuit

.PARAM PI = 3.14159265359
.PARAM heartperiod = <<cycle>>
.PARAM activepeaktime  = <<timetopeaktension>>
.PARAM freq1 = 1 / heartperiod
.PARAM freq2 = 2 / heartperiod
.PARAM freq3 = 3 / heartperiod
.PARAM freq4 = 4 / heartperiod
.PARAM trackrelaxphase = 0
.PARAM lvregurgitation = <<lvregurger>>
.PARAM lvregurgitationvalveratio = <<lvregurgevalveratio>>
.PARAM rvregurgitation = <<rvregurger>>
.PARAM rvregurgitationvalveratio = <<rvregurgevalveratio>>

.func manmod(shorttime) {shorttime - floor(shorttime / heartperiod) * heartperiod}
.func disfrompeak(xtime,peaktime,width) {min( abs( manmod(xtime) - peaktime) , heartperiod - abs( manmod(xtime) - peaktime))}
.func cossq(xtime,amp,peaktime,width) {amp * cos( PI * disfrompeak( xtime , peaktime , width ) / width)^2}

.model valve sidiode(Roff=10k Ron=1m Rrev=10 Vfwd=0.1 Vrev=1k Revepsilon=0.2 Epsilon=0.2)

.subckt vein in out rval=100k lval=1n
R1 1  out    r = rval
L1 in 1    l = lval
.ends vein

Vlaprobe lagnd lagnd2 dc 0
Vraprobe ragnd ragnd2 dc 0
Vlvprobe lv    lvgnd  dc 0
Vrvprobe rvgnd rvgnd2 dc 0

Irvu1   rv       rvgnd   SIN(0 <<rvuamp1>> freq1 0 0 <<rvuphase1>>)
*Irvu2   rv       rvgnd   SIN(0 <<rvuamp2>> freq2 0 0 <<rvuphase2>>)
*Irvu3   rv       rvgnd   SIN(0 <<rvuamp3>> freq3 0 0 <<rvuphase3>>)
*Irvu4   rv       rvgnd   SIN(0 <<rvuamp4>> freq4 0 0 <<rvuphase4>>)

Cra    ra       ragnd   <<rac>> 
Cla    la       lagnd   <<lac>> 

alvu1 %v[lvgenerator] pwl_input
.model pwl_input filesource (file="<<lvufile>>" amploffset=[0] amplscale=[1] timeoffset=0 timescale=1 timerelative=false amplstep=false)

*Blvu2  lvgenerator gnd V = v(lvgenerator0) + v(lvgenerator1)
*alvu20 gnd lvvol %v(lvgenerator0) lvutabmod0
*.model lvutabmod0 table2d (offset=0.0 gain=1 order=3 file="<<lvutablebasefile>>")
*alvu21 lvvol timecyclic %v(lvgenerator1) lvutabmod
*alvu22 lvvol phasetime %v(lvgenerator1) lvutabmod
*.model lvutabmod table2d (offset=0.0 gain=1 order=3 file="<<lvutablefile>>")

.if (trackrelaxphase == 1)
Bestphase lvestphase gnd V = v(timecyclic)/activepeaktime
Blvrisecurrent gnd lvcurrentphase I =  ((v(timecyclic) <= activepeaktime) ? (v(lvcurrentphase) >= (1 - (3 * <<stepTime>> * v(lvrisetemp)))  ? (1-v(lvcurrentphase))/(3 * <<stepTime>> * v(lvrisetemp))*v(lvrisetemp) : v(lvrisetemp) ) : 0)
Blvrisetemp lvrisetemp gnd V = 1/activepeaktime*10
Blvfallcurrent lvcurrentphase gnd I = (v(timecyclic) < activepeaktime) ? 0 : v(lvfalltemp)
Blvfalltemp lvfalltemp gnd V =  1/v(lvtr)

alvpressgrad  lvcurrentphase gnd lvtrcap
.model lvtrcap capacitor (c=1 ic=0)
alvtr gnd lvvol %v(lvtr) lvutabtrmod
.model lvutabtrmod table2d (offset=0.0 gain=1 order=3 file="<<lvtrtablefile>>")
Blvphase lvphase gnd V = max(0,min(1,v(lvcurrentphase)))
Btime2 phasetime gnd V =  (v(timecyclic) > activepeaktime) ? (activepeaktime + v(lvtr) * (1-v(lvcurrentphase))) : v(timecyclic)

.else
Vpassphasetime phasetime timecyclic dc 0
.endif

Etime timecyclic gnd vol = 'manmod(TIME)'

Blavol  lavol gnd I = -i(Vlaprobe) 
alavolconvert  lavol gnd lavolconvertcap
.model lavolconvertcap capacitor (c=1 ic=<<lainitvol>>)

Bravol  ravol gnd I = -i(Vraprobe) 
aravolconvert  ravol gnd ravolconvertcap
.model ravolconvertcap capacitor (c=1 ic=<<rainitvol>>)

Blvvol  lvvol gnd I = -i(Vlvprobe) 
alvvolconvert  lvvol gnd lvvolconvertcap
.model lvvolconvertcap capacitor (c=1 ic=<<lvinitvol>>)

Brvvol  rvvol gnd I = -i(Vrvprobe) 
arvvolconvert  rvvol gnd rvvolconvertcap
.model rvvolconvertcap capacitor (c=1 ic=<<rvinitvol>>)

Blvu   lvgnd   lvgnd2  <<lvinputvar>> = v(lvgenerator)
Vlvu   lvgnd2   gnd  dc 0
*Elvu   lvgnd2  gnd     vol = 'v(lv)'
Ervu   rvgnd2  gnd     vol = 'v(rv)'

Elau   lagnd2  gnd     vol = 'cossq( TIME ,<<laamp>>,<<lapeaktime>>,<<lawidth>>)'
Erau   ragnd2  gnd     vol = 'cossq( TIME ,<<raamp>>,<<rapeaktime>>,<<rawidth>>)'

Xlalavalv  la  lavalvp1    vein  rval=<<lalavalvr>>    lval=<<lalavalvl>>
Vlalavalv  lavalvp1 lavalvp2 dc 0
Blalavalv  lavalvp2 lavalv V=' <<lalavalvk>> * ( i(Vlalavalv) ^2 )^( <<lalavalvb>> / 2) * sgn( i(Vlalavalv) ) '
Xlvlvvalv  lv  lvvalvp1    vein  rval=<<lvlvvalvr>>    lval=<<lvlvvalvl>>
Vlvlvvalv  lvvalvp1 lvvalvp2 dc 0
Blvlvvalv  lvvalvp2 lvvalv V=' <<lvlvvalvk>> * ( i(Vlvlvvalv) ^2 )^( <<lvlvvalvb>> / 2) * sgn( i(Vlvlvvalv) ) '
Xraravalv  ra  ravalvp1    vein  rval=<<raravalvr>>    lval=<<raravalvl>>
Vraravalv  ravalvp1 ravalvp2 dc 0
Braravalv  ravalvp2 ravalv V=' <<raravalvk>> * ( i(Vraravalv) ^2 )^( <<raravalvb>> / 2) * sgn( i(Vraravalv) ) '
Xrvrvvalv  rv  rvvalvp1    vein  rval=<<rvrvvalvr>>    lval=<<rvrvvalvl>>
Vrvrvvalv  rvvalvp1 rvvalvp2 dc 0
Brvrvvalv  rvvalvp2 rvvalv V=' <<rvrvvalvk>> * ( i(Vrvrvvalv) ^2 )^( <<rvrvvalvb>> / 2) * sgn( i(Vrvrvvalv) ) '


alv   lvvalv   aa    valve
.if (lvregurgitation > 0)
Rlvregurgitation lv lvregurp1             r = lvregurgitation
Vlvregurgitation lvregurp1 lavalvp1       dc 0
.elseif (lvregurgitationvalveratio > 0)
Vlvregurgitation  lv          lvregurp1   dc 0
Blvregurgitation  lvregurp1   lvregurp2   V=' <<lalavalvk>> / lvregurgitationvalveratio * ( i(Vlvregurgitation) ^2 )^( <<lalavalvb>> / 2) * sgn( i(Vlvregurgitation) ) '
alvregurgitation  lvregurp2   lavalvp1    valve
.else
Vlvregurgitation  lvregurp1   gnd         dc 0
.endif
ala   lavalv   lv    valve
arv   rvvalv   pa1   valve
.if (rvregurgitation > 0)
Rrvregurgitation rv rvregurp1             r = rvregurgitation
Vrvregurgitation rvregurp1                rvvalvp1 dc 0
.elseif (rvregurgitationvalveratio > 0)
Vrvregurgitation  rv          rvregurp1   dc 0
Brvregurgitation  rvregurp1   rvregurp2   V=' <<raravalvk>> / rvregurgitationvalveratio * ( i(Vrvregurgitation) ^2 )^( <<raravalvb>> / 2) * sgn( i(Vrvregurgitation) ) '
arvregurgitation  rvregurp2   ravalvp1    valve
.else
Vrvregurgitation  rvregurp1   gnd         dc 0
.endif
ara   ravalv   rv    valve
afo   fovalv   la    valve

Caa   aa    gnd    <<aac>>    
Cao1  ao1   gnd    <<ao1c>>   
Cao2  ao2   gnd    <<ao2c>>   
Cao3  ao3   gnd    <<ao3c>>   
Cao4  ao4   gnd    <<ao4c>>   
Cbr   br    gnd    <<brc>>    
Cca   ca    gnd    <<cac>>    
Cub   ub    gnd    <<ubc>>    
Che   he    gnd    <<hec>>    
Cinte inte  gnd    <<intec>> 
Civc  ivc   gnd    <<ivcc>>   
Ckid  kid   gnd    <<kidc>>  
Cleg  leg   gnd    <<legc>>   
Clung lung  gnd    <<lungc>>  
Cpa1  pa1   gnd    <<pa1c>>   
Cpa2  pa2   gnd    <<pa2c>>   
Cplac plac  gnd    <<placc>>  
Csvc  svc   gnd    <<svcc>>  
Cuv   uv    gnd    <<uvc>>   

Xcabr     ca    br     vein  rval=<<cabrr>>     lval=<<cabrl>>
Xbrsvc    br    svc    vein  rval=<<brsvcr>>    lval=<<brsvcl>>
Xubsvc    ub    svc    vein  rval=<<ubsvcr>>    lval=<<ubsvcl>>
Xao1ca    ao1   ca     vein  rval=<<ao1car>>    lval=<<ao1cal>>
Xao1ub    ao1   ub     vein  rval=<<ao1ubr>>    lval=<<ao1ubl>>
Xsvcra    svc   ra     vein  rval=<<svcrar>>    lval=<<svcral>>
Xpa1pa2   pa1   pa2    vein  rval=<<pa1pa2r>>   lval=<<pa1pa2l>>
Xpa2lung  pa2   lung   vein  rval=<<pa2lungr>>  lval=<<pa2lungl>>
Xlungla   lung  la     vein  rval=<<lunglar>>   lval=<<lunglal>>
Xaaao1    aa    ao1    vein  rval=<<aaao1r>>    lval=<<aaao1l>>
Xao1ao2   ao1   ao2    vein  rval=<<ao1ao2r>>   lval=<<ao1ao2l>>
Xao2ao3   ao2   ao3    vein  rval=<<ao2ao3r>>   lval=<<ao2ao3l>>
Xao3ao4   ao3   ao4    vein  rval=<<ao3ao4r>>   lval=<<ao3ao4l>>
Xao3kid   ao3   kid    vein  rval=<<ao3kidr>>   lval=<<ao3kidl>>
Xao3he    ao3   he     vein  rval=<<ao3her>>    lval=<<ao3hel>>
Xao3inte  ao3   inte   vein  rval=<<ao3inter>>  lval=<<ao3intel>>
Xao4leg   ao4   leg    vein  rval=<<ao4legr>>   lval=<<ao4legl>>
Xao4plac  ao4   plac   vein  rval=<<ao4placr>>  lval=<<ao4placl>>
Xkidivc   kid   ivc    vein  rval=<<kidivcr>>   lval=<<kidivcl>>
Xintehe   inte  he     vein  rval=<<inteher>>   lval=<<intehel>>
Xlegivc   leg   ivc    vein  rval=<<legivcr>>   lval=<<legivcl>>
Xplacuv   plac  uv     vein  rval=<<placuvr>>   lval=<<placuvl>>
Xuvhe     uv    he     vein  rval=<<uvher>>     lval=<<uvhel>>
Xheivc    he    ivc    vein  rval=<<heivcr>>    lval=<<heivcl>>
Xivcra    ivc   ra     vein  rval=<<ivcrar>>    lval=<<ivcral>>

Xda       pa2   ao2p1    vein  rval=<<dar>>    lval=<<dal>>
Vda  ao2p1 ao2p2 dc 0
Bda  ao2p2 ao2 V=' <<dak>> * ( i(Vda) ^2 )^( <<dab>> / 2) * sgn( i(Vda) ) '
Xdv       uv    ivcp1    vein  rval=<<dvr>>    lval=<<dvl>>
Vdv  ivcp1 ivcp2 dc 0
Bdv  ivcp2 ivc V=' <<dvk>> * ( i(Vdv) ^2 )^( <<dvb>> / 2) * sgn( i(Vdv) ) '
Xfo       ivc   fovalvp1 vein  rval=<<for>>    lval=<<fol>>
Vfo  fovalvp1 fovalvp2 dc 0
Bfo  fovalvp2 fovalv V=' <<fok>> * ( i(Vfo) ^2 )^( <<fob>> / 2) * sgn( i(Vfo) ) '

.options savecurrents

.ic v(la)= <<vla0>> v(ra)= <<vra0>>
.tran <<stepTime>> <<stopTime>>
*.print tran v(lv) i(Vlvprobe)


.control
set controlswait
set filetype=ascii
set wr_vecnames
run
wrdata <<outfile>> v(lv) v(lvvol) v(la) v(rv) v(ra) v(pa1) v(aa) i(Vlvprobe) v(phasetime)
.endc 
.end
